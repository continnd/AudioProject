module AudioRecorder(
  // Clock Input (50 MHz)
  input CLOCK_50, // 50 MHz
  input CLOCK_27, // 27 MHz
  //  Push Buttons
  input  [3:0]  KEY,
  //  DPDT Switches 
  input  [17:1]  SW,
  //  7-SEG Displays
  // TV Decoder
  output TD_RESET, // TV Decoder Reset
  // I2C
  inout  I2C_SDAT, // I2C Data
  output I2C_SCLK, // I2C Clock
  // Audio CODEC
  output/*inout*/ AUD_ADCLRCK, // Audio CODEC ADC LR Clock
  input	 AUD_ADCDAT,  // Audio CODEC ADC Data
  output /*inout*/  AUD_DACLRCK, // Audio CODEC DAC LR Clock
  output AUD_DACDAT,  // Audio CODEC DAC Data
  inout	 AUD_BCLK,    // Audio CODEC Bit-Stream Clock
  output AUD_XCK,     // Audio CODEC Chip Clock
  inout [15:0]SRAM_DQ,
  output reg [17:0]SRAM_ADDR,
  output SRAM_WE_N,
  output SRAM_UB_N,
  output SRAM_LB_N,
  output SRAM_CE_N,
  output SRAM_OE_N,
  input rst
);

reg[15:0] mem_in;
wire [6:0] myclock;
wire RST;
assign RST = KEY[0];

assign SRAM_DQ = 16'hzzzz;
assign SRAM_UB_N = 1'b0;
assign SRAM_LB_N = 1'b0;
assign SRAM_CE_N = 1'b0;
assign SRAM_OE_N = 1'b0;

// reset delay gives some time for peripherals to initialize
wire DLY_RST;
Reset_Delay r0(	.iCLK(CLOCK_50),.oRESET(DLY_RST) );

assign	TD_RESET = 1'b1;  // Enable 27 MHz

VGA_Audio_PLL 	p1 (	
	.areset(~DLY_RST),
	.inclk0(CLOCK_27),
	.c0(VGA_CTRL_CLK),
	.c1(AUD_CTRL_CLK),
	.c2(VGA_CLK)
);

I2C_AV_Config u3(	
//	Host Side
  .iCLK(CLOCK_50),
  .iRST_N(KEY[0]),
//	I2C Side
  .I2C_SCLK(I2C_SCLK),
  .I2C_SDAT(I2C_SDAT)	
);

assign	AUD_ADCLRCK	=	AUD_DACLRCK;
assign	AUD_XCK		=	AUD_CTRL_CLK;

audio_clock u4(	
//	Audio Side
   .oAUD_BCK(AUD_BCLK),
   .oAUD_LRCK(AUD_DACLRCK),
//	Control Signals
  .iCLK_18_4(AUD_CTRL_CLK),
   .iRST_N(DLY_RST)	
);

wire [15:0] audio_inL, audio_inR;
reg [15:0] audio_outL,audio_outR;

always @(posedge AUD_DACLRCK)
begin
	if(!SW[17])
	begin
		audioR <= audio_inR;
		mem_in <= audio_inR;
		
		if(!rst)
		begin
			SEL_Addr <= 18'd0;
			counter <= 4'd0;
		end
		else
		begin
				SEL_Addr <= SEL_Addr + 1'b1;
		end
		
	end
	else
	begin
		audioR <= SRAM_DQ;
		
		if(!rst)
		begin
			SEL_Addr <= 1'd0;
		end
		else
		begin
			SEL_Addr <= SEL_Addr + 1'b1;
		end
		
	end
end
always @(negedge AUD_DACLRCK)
begin
	if(!SW[17])
	begin
		audioL <= audio_inL;
	end
	else
	begin
		audioL <= SRAM_DQ;
	end
end

reg [15:0]audioL;
reg [15:0]audioR;
reg [4:0] counter;
reg write;
reg[17:0] SEL_Addr;
	

assign SRAM_DQ = SW[17] ? 16'hzzzz : mem_in;
assign SRAM_ADDR = SEL_Addr;
assign SRAM_WE_N = SW[17];
	
assign audio_outL = audioL;
assign audio_outR = audioR;


audio_converter u5(
	// Audio side
	.AUD_BCK(AUD_BCLK),       // Audio bit clock
	.AUD_LRCK(AUD_DACLRCK), // left-right clock
	.AUD_ADCDAT(AUD_ADCDAT),
	.AUD_DATA(AUD_DACDAT),
	// Controller side
	.iRST_N(DLY_RST),  // reset
	.AUD_outL(audio_outL),
	.AUD_outR(audio_outR),
	.AUD_inL(audio_inL),
	.AUD_inR(audio_inR),
);

endmodule
